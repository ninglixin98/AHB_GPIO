`ifndef RKV_GPIO_ELEMENT_SEQUENCES_SVH
`define RKV_GPIO_ELEMENT_SEQUENCES_SVH


`include "rkv_gpio_base_element_sequence.sv"
`include "rkv_gpio_single_write_seq.sv"
`include "rkv_gpio_single_read_seq.sv"


`endif // RKV_GPIO_ELEMENT_SEQUENCES_SVH
