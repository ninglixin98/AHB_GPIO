`ifndef RKV_GPIO_PKG_SV
`define RKV_GPIO_PKG_SV

package rkv_gpio_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import lvc_ahb_pkg::*;

  `include "rkv_gpio_defines.sv"
  `include "rkv_gpio_reg.sv"
  `include "rkv_gpio_config.sv"
  `include "rkv_gpio_reg_adapter.sv"
  `include "rkv_gpio_subscriber.sv"
  `include "rkv_gpio_cov.sv"
  `include "rkv_gpio_scoreboard.sv"
  `include "rkv_gpio_virtual_sequencer.sv"
  `include "rkv_gpio_env.sv"
  `include "rkv_gpio_seq_lib.svh"
  `include "rkv_gpio_tests.svh"

endpackage



`endif // RKV_GPIO_PKG_SV
